`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/04/2024 01:03:47 PM
// Design Name: 
// Module Name: clock
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module clock(
input enable,
input reset,
input mode,
output [3:0] timer100ms,
output [3:0] timer10ms,
output [3:0] timer1sec,
output [3:0] timer10sec,
output [3:0] timer1min,
output [3:0] timer10min
    );
    
    
    
endmodule

